library ieee;

use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity mm_linear_correction_tb is
  -- generic ();
end entity;

architecture testbench of mm_linear_correction_tb is
begin
end;